library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Lista1Ex1 is
Port(
  a : in STD_LOGIC;	
  b : in STD_LOGIC;
  c : out STD_LOGIC
);
end Lista1Ex1;

architecture Behavioral of Lista1Ex1 is

begin

C <= a or (a and b);

end Behavioral;
